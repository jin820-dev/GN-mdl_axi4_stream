// ------------------------------------------------------------
// File    : util_task.svh
// Author  : jin820
// Created : 2026-01-01
// Updated :
// History:
// 2026-01-01  Initial version
// ------------------------------------------------------------

task automatic test_task();
    $display("Hello World");
endtask
